// file: common_pkg.sv
package common_pkg;
      bit running = 1; // running flag to stop clock 
	  real clk_rx_period = 0.27125;
endpackage : common_pkg
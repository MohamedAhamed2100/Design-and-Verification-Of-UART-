// file: common_pkg.sv
package common_pkg;
      bit running = 1; // running flag to stop clock 
endpackage : common_pkg